module button_test_circuit(
    input clk,
    input reset_n,
    input button_in,
    output [7:0] AN,
    output [6:0] sseg,
    output DP
);

endmodule